module top_module( input in, output out );
//type1//
assign out = ~in;
//type2//
  //not(out,in);
endmodule

