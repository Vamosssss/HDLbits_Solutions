module top_module(
    input [31:0] a,
    input [31:0] b,
    input sub,
    output [31:0] sum
);
    wire cout1, cout2;
    wire [15:0]sum1, sum2;
    wire [31:0] b_xor;
    assign b_xor = {32{sub}}^b;
    
    add16 inst1(
        .a (a[15:0]),
        .b (b_xor[15:0]),
        .cin (sub),
        .cout (cout1),
        .sum (sum1)
    );
    
    add16 inst2(
        .a (a[31:16]),
        .b (b_xor[31:16]),
        .cin (cout1),
        .cout (cout2),
        .sum (sum2)
    );
    
    assign sum = {sum2,sum1};
    
    
endmodule
